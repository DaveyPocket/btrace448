library ieee;
use ieee.std_logic_1164.all;

package pongpack is
	type color_t is (black, red, green, yellow, blue, magenta, cyan, white);
end pongpack;
